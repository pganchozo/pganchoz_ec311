`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:54:00 04/15/2019 
// Design Name: 
// Module Name:    Top 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Top(clk_in, rst, clr, ent, change, led, AN, sw, seven_out);

input clk_in, rst, clr, ent, change;
input [3:0] sw; 

output reg [5:0] led;
output [3:0] AN;
output [6:0] seven_out;



//ASM asm( 

endmodule
